package request_acknowledge_package;

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "request_acknowledge_item.svh"
`include "req_ack_driver.svh"
`include "req_ack_driver_slv.svh"
`include "req_ack_monitor.svh"
`include "req_ack_sequencer.svh"
`include "req_ack_agent.svh"
`include "req_ack_scoreboard.svh"
`include "req_ack_enviroment.svh"
`include "ra_sequence.svh"
`include "ra_sequence_1.svh"
`include "ra_sequence_2.svh"
`include "ra_sequence_3.svh"
`include "req_ack_test.svh"
`include "req_ack_test_1.svh"
`include "req_ack_test_2.svh"


    
endpackage: request_acknowledge_package